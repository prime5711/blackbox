domain localdomain broadcast
